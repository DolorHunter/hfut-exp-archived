library verilog;
use verilog.vl_types.all;
entity CPU_tb is
end CPU_tb;
