library verilog;
use verilog.vl_types.all;
entity PC_tb is
end PC_tb;
