library verilog;
use verilog.vl_types.all;
entity decoder38_tb is
end decoder38_tb;
