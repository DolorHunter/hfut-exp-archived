library verilog;
use verilog.vl_types.all;
entity mux41_tb is
end mux41_tb;
