library verilog;
use verilog.vl_types.all;
entity ALU_tb is
end ALU_tb;
